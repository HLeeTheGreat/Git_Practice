module first();


endmodulel;
